module router_sync(clock,resetn,data_in,detect_add,full_0,full_1,full_2,empty_0,empty_1,empty_2,write_enb_reg,read_enb_0,read_enb_1,read_enb_2,write_enb,fifo_full,vld_out_0,vld_out_1,vld_out_2,soft_reset_0,soft_reset_1,soft_reset_2);


input clock,resetn,detect_add,full_0,full_1,full_2,empty_0,empty_1,empty_2,write_enb_reg,read_enb_0,read_enb_1,read_enb_2;
input [1:0]data_in;
output reg[2:0]write_enb;
output reg fifo_full,soft_reset_0,soft_reset_1,soft_reset_2;
output vld_out_0,vld_out_1,vld_out_2;

//declaring internal variable for internal address storing
  reg [1:0] int_addr_reg;  // afterwards we can use it to generate the write_enb

  //declaring counter identifiers for soft_reset which counts 30 clock cyles delay if no respose than it will be developed
  reg[4:0]count_0,count_1,count_2;
  
   //logic for latching adder
  always@(posedge clock)
  begin
    if(!resetn)
    int_addr_reg<=2'b0;  // as active low reset, written 
    else if(detect_add)
    int_addr_reg<=data_in; // as data_in is wire type
  end


  //-----------------------------------Valid Byte block----------------------------------

assign vld_out_0 = (~empty_0);  //it tells that there is a valid byte available for the destination client nerwork 0
assign vld_out_1 = (~empty_1);
assign vld_out_2 = (~empty_2);

  
//-----------------------------------Soft Reset block----------------------------------
  
  
  
//-----------Address decoding & fifo empty ---------------

/*        
    in the below following case only the fifo_full = 1'b1;
    if internal address if 00 and full_0 = 1 then, fifo_full = 1
    if internal address if 01 and full_1 = 1 then, fifo_full = 1
    if internal address if 10 and full_2 = 1 then, fifo_full = 1
        basically from the above conditions we can say that at a particular internal address fifo_full = fifo_X, X = 0,1,2.
    */ 
always@(*)
  begin
    case(int_addr_reg)  // it is dependent in data_in
      2'b00:begin
	          fifo_full<=full_0;
	          if(write_enb_reg) // this write_enb_reg is generated by the fsm.
	          write_enb<=3'b001;  //it is in book pg.no: 18 where due to data_in the write_enb is detected.
	          else
	          write_enb<=3'b0;
	        end

      2'b01:begin
	          fifo_full<=full_1;
	          if(write_enb_reg)
	          write_enb<=3'b010;
	          else
	          write_enb<=3'b0;
	        end

      2'b10:begin
	          fifo_full<=full_2;
	          if(write_enb_reg)
	          write_enb<=3'b100;
	          else
	          write_enb<=3'b0;
	        end
      default:begin
	          fifo_full<=1'b0;
	          write_enb<=1'b0;
	        end
    endcase
  end
  

//-----------------------------------Soft Reset block----------------------------------

// as we are getting some warnings,description: combinational and sequential parts of fsm, it means we can't use same variable to check the condition and update them in the condition block itself, 
  wire c_0 = (count_0==5'd29) ? 1'b1 : 1'b0;  // instead of using these in the respective 'if' statement condition, we have to assign like this, to avoid the above stated warrning
  wire c_1 = (count_1==5'd29) ? 1'b1 : 1'b0;
  wire c_2 = (count_2==5'd29) ? 1'b1 : 1'b0; 


 // for fifo_0
always@(posedge clock)
  begin
  
  if(!resetn)
  begin
  count_0<=5'b0;
  soft_reset_0<=1'b0;
  end

  else if(vld_out_0)
  begin
  if(!read_enb_0)
   
    begin
    if(count_0==5'd29)   // 30 clock cycles
      begin
      soft_reset_0<=1'b1;
      count_0<=5'b0;
      end
    else
      begin
      soft_reset_0<=1'b0;
      count_0<=count_0+1'b1; // at valid out is high, it is generated based on the empty signal
      end
    end
  else
  count_0<=5'b0;
  end
  end

 // for fifo_1
always@(posedge clock)
  begin
  
  if(!resetn)
  begin
  count_1<=5'b0;
  soft_reset_1<=1'b0;
  end

  else if(vld_out_1)
  begin
  if(!read_enb_1)
   
    begin
    if(c_1)
      begin
      soft_reset_1<=1'b1;
      count_1<=5'b0;
      end
    else
      begin
      soft_reset_1<=1'b0;
      count_1<=count_1 + 1'b1;
      end
    end
  else
  count_1<=5'b0;
  end
  end

 // for fifo_2
always@(posedge clock)
  begin
  
  if(!resetn)
  begin
  count_2<=5'b0;
  soft_reset_2<=1'b0;
  end

  else if(vld_out_2)
  begin
  if(!read_enb_2)
   
    begin
    if(c_2)
      begin
      soft_reset_2<=1'b1;
      count_2<=1'b0;
      end
    else
      begin
      soft_reset_2<=1'b0;
      count_2<=count_2+1'b1;
      end
    end
  else
  count_2<=1'b0;
  end
  end

endmodule



// //************ test bench  at time 45:00 in Q & A *****************/
// `timescale 1ns/1ps
// module router_sync_tb();
// 	wire [2:0]write_enb;
// 	wire fifo_full;
// 	wire vld_out_0,vld_out_1,vld_out_2;
// 	wire soft_reset_0,soft_reset_1,soft_reset_2;
// 	reg  clock,resetn,detect_add;
// 	reg  [1:0]data_in;
// 	reg  full_0,full_1,full_2;
// 	reg  empty_0,empty_1,empty_2;
//         reg write_enb_reg;
//         reg read_enb_0,read_enb_1,read_enb_2;
//         parameter T=20;
    
// router_sync DUT(clock,resetn,data_in,detect_add,full_0,full_1,full_2,empty_0,empty_1,empty_2,write_enb_reg == 1'b1,read_enb_0,read_enb_1,read_enb_2,write_enb,fifo_full,vld_out_0,vld_out_1,vld_out_2,soft_reset_0,soft_reset_1,soft_reset_2);
	
//           initial 
//             begin
//               clock=1'b0;
//               forever #(T/2) clock = ~clock;
//             end      
// //task initialize	
//            task initialize;
//  	        begin
// 		     {detect_add,data_in,full_0,full_1,full_2}=0;
// 		     {write_enb_reg,read_enb_0,read_enb_1,read_enb_2,empty_0,empty_1,empty_2}=0;

// 	        end
// 	       endtask
// //task reset
// 	      task reset_dut();
//                   begin
//                     @(negedge clock)  //because it is an active low reset, specified in the data sheet
//                       resetn=1'b0; 
// 		            @(negedge clock)
//                       resetn=1'b1; 
//                   end
//               endtask
// //task read_enb_X ,here X = 0,1,2
//                 task readenb(input r1,r2,r3);
//                    begin
//                         {read_enb_0,read_enb_1,read_enb_2}={r1,r2,r3};
// 		            end 
//                endtask
// //task input and detect addresee
//                  task input_detect (input [1:0] d1,input detect_ad1);
//                     begin
//                       data_in=d1;
// 		              detect_add=detect_ad1;
//                     end
//       		endtask
// //task fifo_full     
// 		task fifo_ful(input f1,f2,f3);
//                     begin
//                       full_0=f1;
//                       full_1=f2;
//                       full_2=f3;
//                      end
//                 endtask
// //task empty
//                task empty_dut(input e1,e2,e3);
//                   begin
// 		            empty_0=e1;
// 		            empty_1=e2;
//                 empty_2=e3;
// 		  		  end
// 			    endtask 
  
//   //task write enb reg
//                 task write_enable_reg (input l1);
//                     begin
//                     write_enb_reg =l1;

//                     end
//                endtask
//  initial begin
// 		initialize;
// 		reset_dut;
//     #20;
//      $display("-------------------------------------------------------------------------------------");
//     @(negedge clock)
// 		readenb(1,0,0);  // here, read_enb_3 = 1'b1; "read_enb_0, read_enb_1, read_enb_2" 
//         input_detect(2'b00,1);
//            fifo_ful(0,0,0);   //full_0, full_1, full_2
//         write_enable_reg (1);
//            empty_dut(0,0,0);  // so here in this case i was expecting vld_out_0,vld_out_1,vld_out_2 = 1'b1;
//            #20;
//            reset_dut;
//            #20 @(negedge clock) input_detect(2'b10,1);
//            write_enable_reg(1'b1);
//            // here the expected output is write_enb = 3'b100
//         $display("--------------------------------at full_1 then, fifo_full = 1-----------------------------------------------------");
//            // now to verify whether the full signal is generated properly
//            #20 @(negedge clock) input_detect(2'b01,1);
//            full_0 = 1; //in this case, output fifo_full = 1'b0; due to fact that "data_in" is 2'b01 not 2'b00
//            @(negedge clock) full_2 = 1;  //in this case, output fifo_full = 1'b0; due to fact that "data_in" is 2'b01 not 2'b10
//           @(negedge clock) full_1 = 1;    // here fifo_full = 1'b1; as data_ip is 2'b01
        

//     $display("--------------------------------------soft reset = 0-----------------------------------------------");
//     #310; // as 300+40 simulation time has 15 clock cycles so no soft_reset_0  (ie. 15xT = 15x20 = 300) 
//     read_enb_0 = 1'b1;  // the read enable has to be made within the 30 clock cycles or else the soft reset will be triggered.
//     // if delay is 600 simulation time(instead of 300) after, the read_enb_0 becomes 1 then soft_reset will be triggered before read_end_0 so, after read_end_0 changes so again the soft_reset becomes 0
//     //30 clock cycles means 30xT = 30x20 = 600 simulation time
//     $display("----------------------------soft reset = 1 if there is no change in the inputs-----------------------------");
//     // Note : the soft reset will be active and again in another clock pulse it will be de-active
//                 #900;
//            $finish;
//   end

// initial
//      begin
//        $monitor($time,"-data_in = %b, detect_add = %b, write_enb = %b, write_enb_reg == 1'b1 = %b,full_0 = %b,full_1 = %b,full_2 = %b, fifo_full = %b, vld_out_0 = %b, soft_reset_1 = %b,clk = %b ",data_in,detect_add,write_enb,write_enb_reg,full_0,full_1,full_2,fifo_full,vld_out_0,soft_reset_1,clock);
//        $dumpfile("router_sync_tb.vcd");
//        $dumpvars;
	
//      end
// endmodule
  
